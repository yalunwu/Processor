library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity writeBack is
  port (
	clock
  ) ;
end entity ; 